* Extracted by KLayout on : 05/09/2021 15:51

.SUBCKT basic_opamp
M$1 VDD IBIAS1 \$5 VP sky130_fd_pr__pfet_g5v0d10v5 L=500000U W=25000000U
+ AS=5.1832e+12P AD=9.48755e+12P PS=24440000U PD=53990000U
M$2 VDD IBIAS1 \$1 VP sky130_fd_pr__pfet_g5v0d10v5 L=500000U W=25000000U
+ AS=5.1832e+12P AD=8.6718e+12P PS=24440000U PD=53860000U
M$3 VOUT VB1 \$1 VP sky130_fd_pr__pfet_g5v0d10v5 L=500000U W=10000000U
+ AS=1.8832e+12P AD=3.2673e+12P PS=9440000U PD=23680000U
M$4 IBIAS1 IBIAS1 VDD VP sky130_fd_pr__pfet_g5v0d10v5 L=500000U W=5000000U
+ AS=1.55e+12P AD=1.65e+12P PS=10620000U PD=10660000U
M$5 \$11 VB1 \$5 VP sky130_fd_pr__pfet_g5v0d10v5 L=500000U W=10000000U
+ AS=1.8832e+12P AD=3.4488e+12P PS=9440000U PD=23740000U
M$6 \$5 IBIAS1 IBIAS1 VNB$1 sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=5000000U
+ AS=1.45e+12P AD=1.45e+12P PS=10580000U PD=10580000U
M$7 VOUT VB2 \$9 VNB$1 sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=2500000U
+ AS=725000000000P AD=725000000000P PS=5580000U PD=5580000U
M$8 IBIAS2 IN_pos \$1 VNB$1 sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=25000000U
+ AS=5.1832e+12P AD=7.8948e+12P PS=24440000U PD=53820000U
M$9 GND \$11 \$9 VNB$1 sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=2500000U
+ AS=725000000000P AD=725000000000P PS=5580000U PD=5580000U
M$10 \$8 \$11 GND VNB$1 sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=2500000U
+ AS=725000000000P AD=725000000000P PS=5580000U PD=5580000U
M$11 IBIAS1 IBIAS1 \$1 VNB$1 sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=5000000U
+ AS=1.55e+12P AD=1.5e+12P PS=10620000U PD=10600000U
M$12 \$8 VB2 \$11 VNB$1 sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=2500000U
+ AS=725000000000P AD=725000000000P PS=5580000U PD=5580000U
M$13 IBIAS2 IN_neg \$5 VNB$1 sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=25000000U
+ AS=5.1832e+12P AD=9.4068e+12P PS=24440000U PD=54060000U
.ENDS basic_opamp
