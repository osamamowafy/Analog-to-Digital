.subckt df INN INP Ihys VDD VG VNB VOUT
M1 net1 net1 VDD VP sky130_fd_pr__pfet_g5v0d10v5 l=1e+06u w=1e+06u
M2 net10 net1 VDD VP sky130_fd_pr__pfet_g5v0d10v5 l=1e+06u w=1e+06u
M3 net1 INN net2 VNB sky130_fd_pr__nfet_g5v0d10v5 l=500000u w=1e+06u 
M4 net10 INP net2 VNB sky130_fd_pr__nfet_g5v0d10v5 l=500000u w=1e+06u 
M5 net2 VDD GND VNB sky130_fd_pr__nfet_g5v0d10v5 l=1e+06u  w=500000u
M6 net1 VG net3 VNB sky130_fd_pr__nfet_g5v0d10v5 l=500000u w=2e+06u  
M7 net3 Ihys GND VNB sky130_fd_pr__nfet_g5v0d10v5 l=500000u w=500000u
M8 net10 net8 net3 VNB sky130_fd_pr__nfet_g5v0d10v5 l=500000u w=2e+06u
M18 Ihys Ihys GND VNB sky130_fd_pr__nfet_g5v0d10v5 l=500000u w=500000u

M12 VG net8 VDD VP sky130_fd_pr__pfet_g5v0d10v5 l=500000u w=4e+06u 
M10 net8 net10 VDD VP sky130_fd_pr__pfet_g5v0d10v5 l=500000u w=6e+06u 
M16 VOUT VG VDD VP sky130_fd_pr__pfet_g5v0d10v5 l=500000u w=4e+06u 
M22 VG EN VDD VP sky130_fd_pr__pfet_g5v0d10v5 l=500000u w=4e+06u 
M20 VOUT VG GND VNB sky130_fd_pr__nfet_g5v0d10v5 l=500000u w=2e+06u 
M17 net5 EN GND VNB sky130_fd_pr__nfet_g5v0d10v5 l=500000u w=2e+06u
M13 VG net8 net5 VNB sky130_fd_pr__nfet_g5v0d10v5 l=500000u w=2e+06u 
M11 net8 VDD GND VNB sky130_fd_pr__nfet_g5v0d10v5 l=500000u w=500000u 
.ends

