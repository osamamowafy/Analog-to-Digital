* Extracted by KLayout on : 29/08/2021 23:51

.SUBCKT df
M$1 \$8 \$5 VDD VP sky130_fd_pr__pfet_g5v0d10v5 L=500000U W=6000000U
+ AS=1.74e+12P AD=1.74e+12P PS=12580000U PD=12580000U
M$2 \$3 EN VDD VP sky130_fd_pr__pfet_g5v0d10v5 L=500000U W=4000000U
+ AS=1.16e+12P AD=1.16e+12P PS=8580000U PD=8580000U
M$3 VDD \$8 \$3 VP sky130_fd_pr__pfet_g5v0d10v5 L=500000U W=4000000U
+ AS=1.16e+12P AD=1.16e+12P PS=8580000U PD=8580000U
M$4 \$2 \$2 VDD VP sky130_fd_pr__pfet_g5v0d10v5 L=1000000U W=1000000U
+ AS=290000000000P AD=675000000000P PS=2580000U PD=2350000U
M$5 VDD \$2 \$5 VP sky130_fd_pr__pfet_g5v0d10v5 L=1000000U W=1000000U
+ AS=675000000000P AD=290000000000P PS=2350000U PD=2580000U
M$6 VDD \$3 VOUT VP sky130_fd_pr__pfet_g5v0d10v5 L=500000U W=4000000U
+ AS=1.16e+12P AD=1.16e+12P PS=8580000U PD=8580000U
M$7 \$6 INP \$5 VNB sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=1000000U
+ AS=290000000000P AD=290000000000P PS=2580000U PD=2580000U
M$8 \$2 INN \$6 VNB sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=1000000U
+ AS=290000000000P AD=290000000000P PS=2580000U PD=2580000U
M$9 GND \$3 VOUT VNB sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=2000000U
+ AS=580000000000P AD=580000000000P PS=4580000U PD=4580000U
M$10 \$2 \$3 \$4 VNB sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=2000000U
+ AS=580000000000P AD=580000000000P PS=4580000U PD=4580000U
M$11 \$4 \$8 \$5 VNB sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=2000000U
+ AS=590000000000P AD=570000000000P PS=4590000U PD=4570000U
M$12 \$6 VDD GND VNB sky130_fd_pr__nfet_g5v0d10v5 L=1000000U W=500000U
+ AS=147500000000P AD=72500000000P PS=1590000U PD=790000U
M$13 GND Ihys \$4 VNB sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=500000U
+ AS=72500000000P AD=145000000000P PS=790000U PD=1580000U
M$14 GND Ihys Ihys VNB sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=500000U
+ AS=145000000000P AD=145000000000P PS=1580000U PD=1580000U
M$15 \$8 VDD GND VNB sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=500000U
+ AS=145000000000P AD=145000000000P PS=1580000U PD=1580000U
M$16 \$3 \$8 \$9 VNB sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=2000000U
+ AS=580000000000P AD=580000000000P PS=4580000U PD=4580000U
M$17 \$9 EN GND VNB sky130_fd_pr__nfet_g5v0d10v5 L=500000U W=2000000U
+ AS=580000000000P AD=580000000000P PS=4580000U PD=4580000U
.ENDS df
